* NGSPICE file created from inv_layout.ext - technology: sky130A

.subckt inv_layout
X0 vout vin vss vss sky130_fd_pr__nfet_01v8 ad=0.35 pd=2.7 as=0.35 ps=2.7 w=1 l=0.15
X1 vout vin vdd vdd sky130_fd_pr__pfet_01v8 ad=1.225 pd=7.7 as=1.225 ps=7.7 w=3.5 l=0.15
C0 vin vout 0.11434f
C1 vdd vout 0.36189f
C2 vdd vin 0.17136f
C3 vout vss 0.39129f
C4 vin vss 0.39015f
C5 vdd vss 1.52782f
.ends

