magic
tech sky130A
timestamp 1766481275
<< nwell >>
rect -90 -95 135 355
<< nmos >>
rect 15 -270 30 -170
<< pmos >>
rect 15 -75 30 275
<< ndiff >>
rect -20 -180 15 -170
rect -20 -260 -15 -180
rect 5 -260 15 -180
rect -20 -270 15 -260
rect 30 -180 65 -170
rect 30 -260 40 -180
rect 60 -260 65 -180
rect 30 -270 65 -260
<< pdiff >>
rect -20 260 15 275
rect -20 -60 -15 260
rect 5 -60 15 260
rect -20 -75 15 -60
rect 30 260 65 275
rect 30 -60 40 260
rect 60 -60 65 260
rect 30 -75 65 -60
<< ndiffc >>
rect -15 -260 5 -180
rect 40 -260 60 -180
<< pdiffc >>
rect -15 -60 5 260
rect 40 -60 60 260
<< psubdiff >>
rect -60 -305 105 -300
rect -60 -325 -15 -305
rect 5 -325 40 -305
rect 60 -325 105 -305
rect -60 -330 105 -325
<< nsubdiff >>
rect -60 330 105 335
rect -60 310 -15 330
rect 5 310 40 330
rect 60 310 105 330
rect -60 305 105 310
<< psubdiffcont >>
rect -15 -325 5 -305
rect 40 -325 60 -305
<< nsubdiffcont >>
rect -15 310 5 330
rect 40 310 60 330
<< poly >>
rect 15 275 30 295
rect 15 -110 30 -75
rect -20 -120 30 -110
rect -20 -140 -10 -120
rect 10 -140 30 -120
rect -20 -150 30 -140
rect 15 -170 30 -150
rect 15 -290 30 -270
<< polycont >>
rect -10 -140 10 -120
<< locali >>
rect -60 330 105 335
rect -60 310 -15 330
rect 5 310 10 330
rect 35 310 40 330
rect 60 310 105 330
rect -60 305 105 310
rect -15 275 5 305
rect -20 260 10 275
rect -20 -60 -15 260
rect 5 -60 10 260
rect -20 -75 10 -60
rect 35 260 65 275
rect 35 -60 40 260
rect 60 -60 65 260
rect 35 -75 65 -60
rect 40 -110 60 -75
rect -20 -120 15 -110
rect -20 -140 -10 -120
rect 10 -140 15 -120
rect -20 -150 15 -140
rect 40 -120 90 -110
rect 40 -140 65 -120
rect 85 -140 90 -120
rect 40 -150 90 -140
rect 40 -170 60 -150
rect -20 -180 10 -170
rect -20 -260 -15 -180
rect 5 -260 10 -180
rect -20 -270 10 -260
rect 35 -180 65 -170
rect 35 -260 40 -180
rect 60 -260 65 -180
rect 35 -270 65 -260
rect -15 -300 5 -270
rect -60 -305 105 -300
rect -60 -325 -15 -305
rect 5 -325 10 -305
rect 35 -325 40 -305
rect 60 -325 105 -305
rect -60 -330 105 -325
<< viali >>
rect 10 310 35 330
rect -10 -140 10 -120
rect 65 -140 85 -120
rect 10 -325 35 -305
<< metal1 >>
rect -120 330 165 335
rect -120 310 10 330
rect 35 310 165 330
rect -120 305 165 310
rect -120 -120 15 -110
rect -120 -140 -10 -120
rect 10 -140 15 -120
rect -120 -150 15 -140
rect 55 -120 165 -110
rect 55 -140 65 -120
rect 85 -140 165 -120
rect 55 -150 165 -140
rect -120 -305 165 -300
rect -120 -325 10 -305
rect 35 -325 165 -305
rect -120 -330 165 -325
<< labels >>
rlabel metal1 145 320 145 320 1 vdd
rlabel metal1 145 -315 145 -315 1 vss
rlabel metal1 155 -150 165 -110 1 vout
rlabel metal1 -120 -150 -110 -110 1 vin
<< end >>
